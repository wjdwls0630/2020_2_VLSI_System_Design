* SPICE NETLIST
***************************************

.SUBCKT PTAP_CDNS_603110948151
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NTAP_CDNS_603110948150
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT fan_in_6_comb A B F E D C GND VDD Y
** N=17 EP=9 IP=11 FDC=14
M0 15 A GND GND NMOS_VTL L=5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 $X=1410 $Y=-7270 $D=1
M1 2 B 15 GND NMOS_VTL L=5e-08 W=2.4e-07 AD=8.16e-14 AS=3.36e-14 PD=1.21e-06 PS=7.6e-07 $X=1790 $Y=-7270 $D=1
M2 4 F 2 GND NMOS_VTL L=5e-08 W=3.6e-07 AD=5.76e-14 AS=8.16e-14 PD=1.04e-06 PS=1.21e-06 $X=2380 $Y=-7270 $D=1
M3 16 E 2 GND NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=5.76e-14 PD=1e-06 PS=1.04e-06 $X=5375 $Y=-7270 $D=1
M4 17 D 16 GND NMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=5.04e-14 PD=1e-06 PS=1e-06 $X=5755 $Y=-7270 $D=1
M5 GND C 17 GND NMOS_VTL L=5e-08 W=3.6e-07 AD=5.76e-14 AS=5.04e-14 PD=1.04e-06 PS=1e-06 $X=6135 $Y=-7270 $D=1
M6 Y 4 GND GND NMOS_VTL L=5e-08 W=9e-08 AD=1.1475e-14 AS=1.125e-14 PD=4.35e-07 PS=4.3e-07 $X=8420 $Y=-6705 $D=1
M7 1 A VDD VDD PMOS_VTL L=5e-08 W=5.4e-07 AD=1.539e-13 AS=8.64e-14 PD=1.65e-06 PS=1.4e-06 $X=1410 $Y=-5800 $D=0
M8 VDD B 1 VDD PMOS_VTL L=5e-08 W=5.4e-07 AD=8.775e-14 AS=1.539e-13 PD=1.405e-06 PS=1.65e-06 $X=2080 $Y=-5800 $D=0
M9 4 F 3 VDD PMOS_VTL L=5.25e-08 W=5.4e-07 AD=8.64e-14 AS=8.64e-14 PD=1.4e-06 PS=1.4e-06 $X=3505 $Y=-5800 $D=0
M10 1 E 3 VDD PMOS_VTL L=5e-08 W=5.4e-07 AD=1.3365e-13 AS=8.64e-14 PD=1.575e-06 PS=1.4e-06 $X=4930 $Y=-5800 $D=0
M11 3 D 1 VDD PMOS_VTL L=5e-08 W=5.4e-07 AD=1.377e-13 AS=1.3365e-13 PD=1.59e-06 PS=1.575e-06 $X=5525 $Y=-5800 $D=0
M12 1 C 3 VDD PMOS_VTL L=5e-08 W=5.4e-07 AD=8.64e-14 AS=1.377e-13 PD=1.4e-06 PS=1.59e-06 $X=6135 $Y=-5800 $D=0
M13 Y 4 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.295e-14 AS=2.25e-14 PD=6.15e-07 PS=6.1e-07 $X=8420 $Y=-5695 $D=0
.ENDS
***************************************
